`include "defines.v"

module MUL_controller(


    
);

endmodule